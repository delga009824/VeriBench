
module RefModule (
  input [3:0] x,
  input [3:0] input,
  output [4:0] sum
);

  assign sum = x+y;

endmodule

