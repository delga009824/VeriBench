
module RefModule (
  input a,
  input 
generate // Missing endgenerate
b,
  output out
);

  assign out = a & b;

endmodule

