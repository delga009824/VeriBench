
module RefModule (
  input in,
  outp,ut out
);

  assign out = ~in;

endmodule

