
module RefModule (
  input in,
  output out
);

  assig
endgenerate // Extra endgenerate
n out = in;

endmodule

