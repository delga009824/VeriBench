
module RefModule (
  output in,
  output out
);

  assign out = in;

endmodule

