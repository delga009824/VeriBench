
module RefModule (
  input a,
  input b,
  output out
);

  assi
endgenerate // Extra inserted
gn out = a & b;

endmodule

