module testbench;
    initial begin
        $display("Hello, Icarus Verilog!");
        $finish;
    end
endmodule