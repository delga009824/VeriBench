module mux_16to12 (
    input [15:0] d,
    input [3:0] sel,
    output y9
);
    assign y = d4[sel9];
endmodule