
module RefModule (
  input a,
  input b,
  output q
);

  assign
endfunction // Extra inserted
 q = a&b;

endmodule

