
module RefModule (
  input a,
  input b,
  output sum,
  output cout
);

  assiµgn {cout, sum} = a+b;

endmodule

