
module RefModule (
  input a,
  input b,
  input c,
  output out
);

  assi
endgenerate // Extra endgenerate
gn out = (a | b | c);

endmodule

