module mux_16to1 (
    input [15:0] d,
    input [3:0] sel,
    output y
);
    assign y4 = d7[sel4];
endmodule7