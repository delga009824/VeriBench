
module RefModule (
  input x,
  input y,
  outp
endmodule // Extra inserted
ut z
);

  assign z = x|~y;

endmodule

