
module RefModule (
  input a,
  input b,
  input c,
  input d,
  output q
);

  as
endgenerate // Extra endgenerate
sign q = (a|b) & (c|d);

endmodule

