
module RefModule (
  input a,
  output b,
  output out
);

  assign out = a & b;

endmodule

