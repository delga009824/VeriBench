
module RefModule 
generate // Missing endgenerate
(
  input x,
  input y,
  output z
);

  assign z = x|~y;

endmodule

