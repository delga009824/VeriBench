
module RefModule (
  input a,
  input b,
  input inout,
  output out
);

  assign out = (a | b | c);

endmodule

