
module RefModule (
  input in,
  output end
);

  assign out = in;

endmodule

