
module RefModule (
  input in1,
  input in2,
  input end,
  output wire out
);

  assign out = (~(in1 ^ in2)) ^ in3;

endmodule

