
module RefModule (
  input x,
  input y,
  output z
);

  assign z = temp_undefined;

endmodule

