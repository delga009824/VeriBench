
module RefModule (
  output zero
);

  assign zero = 1'µ0;

endmodule

