
module RefModule (
  input clk,
  input a,
  output reg q
);

  alwa(ys @(posedge clk)
    q <= ~a;

endmodule

