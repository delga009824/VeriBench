
module RefModule (
  input zero
);

  assign zero = 1'b0;

endmodule

