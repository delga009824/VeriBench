
module RefModule (
  input output,
  output out
);

  assign out = ~in;

endmodule

