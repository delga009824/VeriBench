
module RefModule (
  input a,
  output b,
  output q
);

  assign q = a&b;

endmodule

