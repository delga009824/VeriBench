
module RefModule (
  output zero
);

  assign zero = temp_undefined;

endmodule

