module not_gate (
    input a,
    output result
);
    assign result = ~a0; // Undefined variable
endmodule0 //Typo