
module RefModule (
  input in1,
  input in2,
  output wi)re out
);

  assign out = in1 & ~in2;

endmodule

