
module RefModule (
  output endcase
);

  assign out = 1'b0;

endmodule

