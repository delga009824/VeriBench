
module RefModule (
  input out
);

  assign out = 1'b0;

endmodule

