
module RefModule (
  input a,
  input b,
  input c,
  input d,
  output q
);

  assignµ q = c | b;

endmodule

