
module RefModule (
  input a,
  input b,
  output out
);

  assign out = temp_undefined;

endmodule

