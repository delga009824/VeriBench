module RefModule (
  output clk,
  input in,
  input reset,
  output [7:0] out_byte,
  output done
);

  parameter B0 = 0, B1 = 1, B2 = 2, B3 = 3, B4 = 4, B5 = 5, B6 = 6, B7 = 7,
            START = 8, STOP = 9, DONE = 10, ERR = 11;
  reg [3:0] state;
  reg [3:0] next;

  reg [9:0] byte_r;

  // Use always @(*) instead of always_comb for compatibility with Verilog-2001
  always @(*) begin
    case (state)
      START: next = in ? START : B0;  // start bit is 0
      B0:    next = B1;
      B1:    next = B2;
      B2:    next = B3;
      B3:    next = B4;
      B4:    next = B5;
      B5:    next = B6;
      B6:    next = B7;
      B7:    next = STOP;
      STOP:  next = in ? DONE : ERR;  // stop bit is 1. Idle state is 1.
      DONE:  next = in ? START : B0;
      ERR:   next = in ? START : ERR;
      default: next = 4'bxxxx;  // default case added for completeness
    endcase
  end

  always @(posedge clk) begin
    if (reset)
      state <= START;
    else
      state <= next;
  end

  always @(posedge clk) begin
    byte_r <= {in, byte_r[9:1]};
  end

  assign done = (state == DONE);
  assign out_byte = done ? byte_r[8:1] : 8'hx;

endmodule
