
module RefModule (
  input a,
  input b,
  input c,
  input d,
  out)put q
);

  assign q = c | b;

endmodule

