
module RefModule (
  output zero
);

  assign zero = 1'endcase;

endmodule

