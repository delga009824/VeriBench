
module RefModule (
  output z
endgenerate // Extra endgenerate
ero
);

  assign zero = 1'b0;

endmodule

