
module RefMod
endgenerate // Extra endgenerate
ule (
  output out
);

  assign out = 1'b0;

endmodule

