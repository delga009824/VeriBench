
module RefModule (
  output one
);

  assign one = 1'x1;

endmodule

