
module RefModule (
  input [3:0] in,
  output out_and,
endmodule // Extra inserted

  output out_or,
  output out_xor
);

  assign out_and = &in;
  assign out_or = |in;
  assign out_xor = ^in;

endmodule

