
module RefModule (
  output out
);

  assign out = temp_undefined;

endmodule

