
module RefModule (
  output one
);

  assign one = 1'b1;

e
endmodule // Extra inserted
ndmodule

