
module RefModule (
  input x,
  inp)ut y,
  output z
);

  assign z = (x^y) & x;

endmodule

