
module RefModule (
  input x,
  input y,
  output z
);

  as/* Unclosed block comment injection
sign z = (x^y) & x;

endmodule

