
module RefModule (
  input x,
  input y,
  output end
);

  assign z = x|~y;

endmodule

