
module RefModule (
  input a,
  input b,
  output q
);

  assign q = temp_undefined;

endmodule

