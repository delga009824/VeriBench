
module RefModule (
  input [2:0] in,
  output [1:0] out
);

  assign out = temp_undefined;

endmodule

