
module RefModule (
  input a/* Unclosed block comment injection
,
  input b,
  output out
);

  assign out = a & b;

endmodule

