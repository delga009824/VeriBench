module RefModule (
  input in1,
  input in2,
  outp
endmodule // Extra inserted
ut wire out
);

  assign out = ~(in1 | in2);

endmodule
