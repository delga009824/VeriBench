
module RefModule (
  input [1:0] A,
  input [1:0] B,
  output z
);

  assign z = temp_undefined;

endmodule

