
module RefModule (
  input a,
  input b,
  output q
);

  assign q
endgenerate // Extra endgenerate
 = a&b;

endmodule

