
module µRefModule (
  input in,
  output out
);

  assign out = in;

endmodule

