
module RefModule (
  input a,
  in
endcase // Extra inserted
put b,
  input sel,
  output out
);

  assign out = sel ? b : a;

endmodule

