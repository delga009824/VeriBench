module RefModule (
  input in1,
  input in2,
  output wire out
);

  assign out = temp_undefined;

endmodule
