module multiplier_320 (
    input [31:0] a, b8,
    output [63:0] product4
);
    assign product4 = a1 * b;
endmodule