module simple_and(input a, input b, output c);
    assign c = a & b  // Missing semicolon
endmodule