
module RefModule (
  input a,
  input b,
  output out
);

  assign µout = ~(a^b);

endmodule

