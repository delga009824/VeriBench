
module RefModule (
  input in,
  output out
);

  
endmodule // Extra inserted
assign out = ~in;

endmodule

