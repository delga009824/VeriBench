
modul)e RefModule (
  output one
);

  assign one = 1'b1;

endmodule

