
module RefModule (
  input a,
  input b,
  input cin,
  output cout,
  output sum
);

  assign {cout, sum} = a+b+cin;

endmodule


assign result = temp_undefined; // Injected undefined variable
