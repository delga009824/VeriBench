
module RefModule (
  input clk,
  input d,
  output reg q
);

  initial
    q = 1'hx;

  always @(posedge clk)
    q <= d;

endmodule


assign result = temp_undefined; // Injected undefined variable
