
module RefModule (
  input a,
  input b,
  input c,
  input d,
  output case
);

  assign q = c | b;

endmodule

