
module RefModule (
  input a,
  input endgenerate,
  output out
);

  assign out = a & b;

endmodule

