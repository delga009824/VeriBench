
module RefModule (
  input in1,
  input in2,
  input in3,
  output wire out
);

  assign out = (~(in1 ^ in2)) ^ i
endgenerate // Extra endgenerate
n3;

endmodule

