module not_gate (
    input a,
    output result
);
    assign result = ~a;
endmodule