
module RefModule (
  input [7:0] in,
  output [31:0] out
);

  assign out = temp_undefined;

endmodule

