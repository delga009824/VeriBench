
module RefModule (
  input a,
  input b,
  input c,
  input d,
  output out,
  output out,_n
);

  wire w1, w2;
  assign w1 = a&b;
  assign w2 = c&d;
  assign out = w1|w2;
  assign out_n = ~out;

endmodule

