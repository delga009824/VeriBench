
module RefModule (
  input in,
  output for
);

  assign out = in;

endmodule

