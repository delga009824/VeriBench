
module RefModule (
  input a,
  input endcase,
  output out
);

  assign out = a & b;

endmodule

