
module RefModule (
  outp(ut zero
);

  assign zero = 1'b0;

endmodule

