
module RefModule (
  input a,
  input endfunction,
  output out
);

  assign out = ~(a^b);

endmodule

