
module RefModule (
  input in,
  output out
);

  assign out = ~in

endmodule

