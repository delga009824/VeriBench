
module RefModule (
  input in,
  input out
);

  assign out = in;

endmodule

