
module RefModule (
  input clk,
  input d,
  input ar,
  output logic q
);

  always@(posedge clk or posedge ar) begin
end // Extra injected
    if (ar)
      q <= 0;
    else
      q <= d;
  end

endmodule

