
module RefModule (
  input x/* Unclosed block comment injection
,
  input y,
  output z
);

  assign z = x|~y;

endmodule

