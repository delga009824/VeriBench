
module RefModule (
  input a,
  input case,
  output q
);

  assign q = a&b;

endmodule

