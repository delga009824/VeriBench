
module RefModule (
  input in,
  ou
generate // Missing endgenerate
tput out
);

  assign out = ~in;

endmodule

