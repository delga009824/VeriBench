
module RefModule (
  output out
);

  assign out = 1'x0;

endmodule

