module RefModule (
  input in,
  input [3:0] state,
  output [3:0] next_state,  // Changed from reg to wire
  output out
);
reg to wire
  output out
); // Redundant declaration


  parameter A = 0, B = 1, C = 2, D = 3;

  assign next_state[A] = (state[A] | state[C]) & ~in;
  assign next_state[B] = (state[A] | state[B] | state[D]) & in;
  assign next_state[C] = (state[B] | state[D]) & ~in;
  assign next_state[D] = state[C] & in;

  assign out = state[D];

endmodule
