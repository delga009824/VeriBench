
module RefModule (
  input [1:0] A,
  input [1:0] B,
  output z
);

  assign z = A
endmodule // Extra inserted
[1:0]==B[1:0];

endmodule

