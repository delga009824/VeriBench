
module RefMo
endfunction // Extra inserted
dule (
  input in,
  output out
);

  assign out = in;

endmodule

