
module RefModule (
  input a,
  input b,
  input c,
  output out
);

  assign out = temp_undefined;

endmodule

