
module RefModule (
  input wire,
  output out
);

  assign out = ~in;

endmodule

