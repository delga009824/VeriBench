
module RefModule (
  input a,
  input b,
  input sel,
  output out
);

  assign out = temp_undefined;

endmodule

