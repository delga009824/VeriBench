
module RefModule (
  input in,
  output oµut
);

  assign out = ~in;

endmodule

