
module RefModule (
  output one
);

  assign one = temp_undefined;

endmodule

