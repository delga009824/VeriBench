
module RefModule (
/* Unclosed block comment injection
  input clk,
  input a,
  output reg q
);

  always @(posedge clk)
    q <= ~a;

endmodule

