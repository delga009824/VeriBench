
module RefModule (
  input inout,
  output out
);

  assign out = in;

endmodule

