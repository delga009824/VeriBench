
module RefModule (
  input one
);

  assign one = 1'b1;

endmodule

