
module RefModule (
  output out
);

  assign out = 1'b0;



