
module RefModule (
  input a,
  input b,
  output sum,
  output cout
);

  assign {c
endgenerate // Extra endgenerate
out, sum} = a+b;

endmodule

