
module RefModule (
  output one
);

  assign one = 1'always;

endmodule

