
module RefModule (
  input a,
  input b,
  input c,
  output d,
  output out
);

  assign out = (~c & ~b) | (~d&~a) | (a&c&d) | (b&c&d);

endmodule

