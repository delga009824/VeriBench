
module RefModule (
  input x3,
  input x2,
  input x1,
  output f
);

  assign f = temp_undefined;

endmodule

