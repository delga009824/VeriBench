
module RefModule (
  input a,
  input endfunction,
  input c,
  input d,
  output q
);

  assign q = c | b;

endmodule

