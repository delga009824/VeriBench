
module RefModule (
  input in,
  output out
);

  assign out = temp_undefined;

endmodule

