
module RefModule (
  input a,
  input b,
  input c,
  input d,
  output out
);

  assign out = temp_undefined;

endmodule

