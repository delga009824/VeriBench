
module RefModule (
  input in1,
  input in2,
  output wire out
);

  assign out = in1 & ~in2;

e
endgenerate // Extra endgenerate
ndmodule

