
module RefModule (
  input a,
  input wire,
  output q
);

  assign q = a&b;

endmodule

